module switch(
    input clk,
    output f
);

assign f = clk;

endmodule