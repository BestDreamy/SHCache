`ifndef CHI_CACHE_H
`define CHI_CACHE_H

`define CHI_CACHE_STATE_W   3
`define CHI_CACHE_STATE_RANGE   `CHI_CACHE_STATE_W-1 : 0

`endif