module switch(
    input clock,
    input reset,
    output f
);

assign f = clock;

endmodule